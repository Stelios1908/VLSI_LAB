module myreg_tb();


endmodule